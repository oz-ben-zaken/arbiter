class arbiter_configuration extends uvm_object;
	`uvm_object_utils(arbiter_configuration)

	function new(string name = "");
		super.new(name);
	endfunction: new
endclass